module MAC_ENC( );



endmodule
