/* This fifo is modified to support EOD (END OF DATA) signal */
/* EOD indicates packet(frame) end, useful to develop network funciton */

/************************************************************\
 **  Copyright (c) 2011-2021 Anlogic, Inc.
 **  All Right Reserved.
\************************************************************/
/************************************************************\
 ** Log	:	This file is generated by Anlogic IP Generator.
 ** File	:	/home/dudestin/HomemadeSwitch/al_ip/PACKET_FIFO.v
 ** Date	:	2022 07 06
 ** TD version	:	4.4.433
\************************************************************/

`timescale 1ns / 1ps

module PACKET_FIFO (
	rst,
	di, clkw, we,
	do, clkr, re,
	empty_flag, aempty_flag,
	full_flag, afull_flag, 
	// my original signal
	EOD_in, EOD_out
);
	input rst;
	input [7:0] di;
	input clkw, we;
	input clkr,re;

	output [7:0] do;
	output empty_flag, aempty_flag;
	output full_flag, afull_flag;
	// my original signal
	input  wire EOD_in;
	output wire EOD_out;
	
	wire [8:0] new_din;
	wire [8:0] new_dout;

	assign new_din = {di, EOD_in};
	assign do      = new_dout[8:1];
	assign EOD_out = new_dout[0];
	
EG_LOGIC_FIFO #(
 	.DATA_WIDTH_W(9),
	.DATA_WIDTH_R(9),
	.DATA_DEPTH_W(8192),
	.DATA_DEPTH_R(8192),
	.ENDIAN("BIG"),
	.RESETMODE("ASYNC"),
	.E(0),
	.F(8192),
	.ASYNC_RESET_RELEASE("SYNC"),
	.AE(6),
	.AF(6600))
logic_fifo(
	.rst(rst),
	.di(new_din),
	.clkw(clkw),
	.we(we),
	.csw(3'b111),
	.do(new_dout),
	.clkr(clkr),
	.re(re),
	.csr(3'b111),
	.ore(1'b0),
	.empty_flag(empty_flag),
	.aempty_flag(aempty_flag),
	.full_flag(full_flag),
	.afull_flag(afull_flag)

);

endmodule